
module NIOS (
	clk_clk,
	pio_external_export,
	reset_reset_n);	

	input		clk_clk;
	output		pio_external_export;
	input		reset_reset_n;
endmodule
